//------------------------------------------------------------------------------
// fifo_80x2048
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// MIT License
//
// Copyright (c) 2020 homelith
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//------------------------------------------------------------------------------

module fifo_80x2048 (
	input           clk,
	input           xrst,
	input   [79:0]  wdata,
	output          afull,
	output          full,
	input           wval,
	output  [79:0]  rdata,
	output          aempty,
	output          empty,
	input           rval,
	output  [11:0]  usedw
);
	wire    [10:0]  altera_usedw;
	reg             full_1d_r;
	always @ (posedge clk) begin
		full_1d_r <= full;
	end
	assign usedw = {full_1d_r, altera_usedw};
	altera_fifo_80x2048 inst(
		.aclr(~xrst),
		.clock(clk),
		.data(wdata),
		.rdreq(rval),
		.wrreq(wval),
		.almost_empty(aempty),
		.almost_full(afull),
		.empty(empty),
		.full(full),
		.q(rdata),
		.usedw(altera_usedw)
	);
endmodule
